module top ( a , b , c , o);

input a , b , c;

output o;

wire ;

xnor(o,a,b,c);

endmodule
